LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ROM_16 IS 
PORT(
		PC_address: 	IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		INSTRUCTION: 	OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
);
END ROM_16;

ARCHITECTURE ROM_BH OF ROM_16 IS

	CONSTANT instruction0:  STD_LOGIC_VECTOR (15 DOWNTO 0) := "0000000000000001";
	CONSTANT instruction1:  STD_LOGIC_VECTOR (15 DOWNTO 0) := "0000000000000011";
	CONSTANT instruction2:  STD_LOGIC_VECTOR (15 DOWNTO 0) := "0000000000000101";
	CONSTANT instruction3:  STD_LOGIC_VECTOR (15 DOWNTO 0) := "0000000000001001";
	CONSTANT instruction4:  STD_LOGIC_VECTOR (15 DOWNTO 0) := "0000000000100001";
	CONSTANT instruction5:  STD_LOGIC_VECTOR (15 DOWNTO 0) := "0000000001000001";
	CONSTANT instruction6:  STD_LOGIC_VECTOR (15 DOWNTO 0) := "0000000010000001";
	CONSTANT instruction7:  STD_LOGIC_VECTOR (15 DOWNTO 0) := "0000000100000001";
	CONSTANT instruction8:  STD_LOGIC_VECTOR (15 DOWNTO 0) := "0000001000000001";
	CONSTANT instruction9:  STD_LOGIC_VECTOR (15 DOWNTO 0) := "0000010000000001";
	CONSTANT instruction10: STD_LOGIC_VECTOR (15 DOWNTO 0) := "0000100000000001";
	CONSTANT instruction11: STD_LOGIC_VECTOR (15 DOWNTO 0) := "0001000000000001";
	CONSTANT instruction12: STD_LOGIC_VECTOR (15 DOWNTO 0) := "0010000000000001";
	CONSTANT instruction13: STD_LOGIC_VECTOR (15 DOWNTO 0) := "0100000000000001";
	CONSTANT instruction14: STD_LOGIC_VECTOR (15 DOWNTO 0) := "1000000000000001";
	CONSTANT instruction15: STD_LOGIC_VECTOR (15 DOWNTO 0) := "1000000000000011";
	
TYPE ROM_ARRAY IS ARRAY (NATURAL RANGE <>) OF STD_LOGIC_VECTOR (15 DOWNTO 0);
CONSTANT ROM: ROM_ARRAY := (
	instruction0, instruction1, instruction2, instruction3,
	instruction4, instruction5, instruction6, instruction7,
	instruction8, instruction9, instruction10, instruction11,
	instruction12, instruction13, instruction14,instruction15
);

BEGIN 
	PROCESS(PC_address)
	VARIABLE j: integer;
	BEGIN
		j := conv_integer(PC_address);
		INSTRUCTION <= ROM(j);
	END PROCESS;
END ROM_BH;
